library verilog;
use verilog.vl_types.all;
entity mc51_tb is
end mc51_tb;
