//-----------------------------------------------------------------------------------------------------------------------------------------------------------//
//	FILE: 		mc8051_top.v
// 	AUTHOR:		Biggest_apple
// 	
//	ABSTRACT:	
// 	KEYWORDS:	fpga, basic module,signal process
// 
// 	MODIFICATION HISTORY:
//	$Log$
//			Biggest_apple				2024.11.20		Create the project
//-----------------------------------------------------------------------------------------------------------------------------------------------------------//
module mc8051_top(
	input					clk,
	input					reset_n,


);






endmodule