//-----------------------------------------------------------------------------------------------------------------------------------------------------------//
//	FILE: 		basic_periDev.v
// 	AUTHOR:		Biggest_apple
// 	
//	ABSTRACT:	
// 	KEYWORDS:	fpga, basic module,signal process
// 
// 	MODIFICATION HISTORY:
//	$Log$
//			Biggest_apple				2024.12.20		Create the file
//-----------------------------------------------------------------------------------------------------------------------------------------------------------//
`timescale 				1ns/1ps
`include				"global_param.v"
module nvi_periDev(
	input					    clk,
	input					    reset_n,


);


endmodule